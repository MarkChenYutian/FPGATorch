`default_nettype none


module fakemem_readA
  (input logic read, clock, 
   input logic [`ADDR_WIDTH-1:0] address,
   output logic [`BANDWIDTH-1:0][`DATA_WIDTH-1:0] readdata);

  logic [511:0][31:0] mem;

  assign mem[383:0] = {$shortrealtobits(5), $shortrealtobits(2), $shortrealtobits(7), $shortrealtobits(4), $shortrealtobits(1), $shortrealtobits(6), $shortrealtobits(5), $shortrealtobits(7), $shortrealtobits(9), $shortrealtobits(7), $shortrealtobits(4), $shortrealtobits(6), $shortrealtobits(2), $shortrealtobits(10), $shortrealtobits(3), $shortrealtobits(7), $shortrealtobits(10), $shortrealtobits(9), $shortrealtobits(6), $shortrealtobits(5), $shortrealtobits(4), $shortrealtobits(4), $shortrealtobits(5), $shortrealtobits(2), $shortrealtobits(7), $shortrealtobits(8), $shortrealtobits(6), $shortrealtobits(2), $shortrealtobits(9), $shortrealtobits(5), $shortrealtobits(3), $shortrealtobits(4), $shortrealtobits(4), $shortrealtobits(5), $shortrealtobits(3), $shortrealtobits(2), $shortrealtobits(4), $shortrealtobits(7), $shortrealtobits(8), $shortrealtobits(6), $shortrealtobits(6), $shortrealtobits(9), $shortrealtobits(9), $shortrealtobits(10), $shortrealtobits(5), $shortrealtobits(8), $shortrealtobits(1), $shortrealtobits(9), $shortrealtobits(1), $shortrealtobits(6), $shortrealtobits(6), $shortrealtobits(5), $shortrealtobits(8), $shortrealtobits(6), $shortrealtobits(6), $shortrealtobits(2), $shortrealtobits(6), $shortrealtobits(5), $shortrealtobits(5), $shortrealtobits(6), $shortrealtobits(7), $shortrealtobits(9), $shortrealtobits(2), $shortrealtobits(3), $shortrealtobits(5), $shortrealtobits(1), $shortrealtobits(2), $shortrealtobits(1), $shortrealtobits(8), $shortrealtobits(4), $shortrealtobits(4), $shortrealtobits(8), $shortrealtobits(10), $shortrealtobits(3), $shortrealtobits(1), $shortrealtobits(6), $shortrealtobits(6), $shortrealtobits(2), $shortrealtobits(3), $shortrealtobits(8), $shortrealtobits(9), $shortrealtobits(10), $shortrealtobits(5), $shortrealtobits(7), $shortrealtobits(4), $shortrealtobits(10), $shortrealtobits(9), $shortrealtobits(9), $shortrealtobits(2), $shortrealtobits(1), $shortrealtobits(2), $shortrealtobits(5), $shortrealtobits(5), $shortrealtobits(1), $shortrealtobits(8), $shortrealtobits(2), $shortrealtobits(6), $shortrealtobits(3), $shortrealtobits(8), $shortrealtobits(7), $shortrealtobits(3), $shortrealtobits(8), $shortrealtobits(9), $shortrealtobits(10), $shortrealtobits(6), $shortrealtobits(3), $shortrealtobits(8), $shortrealtobits(7), $shortrealtobits(6), $shortrealtobits(7), $shortrealtobits(5), $shortrealtobits(8), $shortrealtobits(9), $shortrealtobits(6), $shortrealtobits(6), $shortrealtobits(10), $shortrealtobits(1), $shortrealtobits(4), $shortrealtobits(1), $shortrealtobits(8), $shortrealtobits(8), $shortrealtobits(8), $shortrealtobits(3), $shortrealtobits(4), $shortrealtobits(5), $shortrealtobits(1), $shortrealtobits(3), $shortrealtobits(10), $shortrealtobits(4), $shortrealtobits(6), $shortrealtobits(2), $shortrealtobits(5), $shortrealtobits(6), $shortrealtobits(2), $shortrealtobits(4), $shortrealtobits(5), $shortrealtobits(5), $shortrealtobits(2), $shortrealtobits(7), $shortrealtobits(8), $shortrealtobits(6), $shortrealtobits(5), $shortrealtobits(4), $shortrealtobits(9), $shortrealtobits(10), $shortrealtobits(1), $shortrealtobits(4), $shortrealtobits(9), $shortrealtobits(1), $shortrealtobits(4), $shortrealtobits(1), $shortrealtobits(4), $shortrealtobits(2), $shortrealtobits(3), $shortrealtobits(10), $shortrealtobits(4), $shortrealtobits(10), $shortrealtobits(5), $shortrealtobits(9), $shortrealtobits(2), $shortrealtobits(4), $shortrealtobits(2), $shortrealtobits(5), $shortrealtobits(3), $shortrealtobits(3), $shortrealtobits(5), $shortrealtobits(5), $shortrealtobits(1), $shortrealtobits(6), $shortrealtobits(10), $shortrealtobits(5), $shortrealtobits(8), $shortrealtobits(1), $shortrealtobits(5), $shortrealtobits(10), $shortrealtobits(3), $shortrealtobits(8), $shortrealtobits(8), $shortrealtobits(5), $shortrealtobits(4), $shortrealtobits(5), $shortrealtobits(10), $shortrealtobits(10), $shortrealtobits(9), $shortrealtobits(7), $shortrealtobits(4), $shortrealtobits(10), $shortrealtobits(3), $shortrealtobits(1), $shortrealtobits(9), $shortrealtobits(6), $shortrealtobits(7), $shortrealtobits(7), $shortrealtobits(10), $shortrealtobits(9), $shortrealtobits(5), $shortrealtobits(3), $shortrealtobits(9), $shortrealtobits(2), $shortrealtobits(9), $shortrealtobits(1), $shortrealtobits(2), $shortrealtobits(4), $shortrealtobits(10), $shortrealtobits(6), $shortrealtobits(2), $shortrealtobits(2), $shortrealtobits(7), $shortrealtobits(6), $shortrealtobits(3), $shortrealtobits(10), $shortrealtobits(1), $shortrealtobits(6), $shortrealtobits(5), $shortrealtobits(1), $shortrealtobits(10), $shortrealtobits(7), $shortrealtobits(1), $shortrealtobits(7), $shortrealtobits(6), $shortrealtobits(3), $shortrealtobits(3), $shortrealtobits(9), $shortrealtobits(5), $shortrealtobits(6), $shortrealtobits(8), $shortrealtobits(5), $shortrealtobits(2), $shortrealtobits(4), $shortrealtobits(6), $shortrealtobits(7), $shortrealtobits(7), $shortrealtobits(9), $shortrealtobits(8), $shortrealtobits(2), $shortrealtobits(1), $shortrealtobits(5), $shortrealtobits(6), $shortrealtobits(3), $shortrealtobits(10), $shortrealtobits(10), $shortrealtobits(2), $shortrealtobits(9), $shortrealtobits(7), $shortrealtobits(5), $shortrealtobits(8), $shortrealtobits(4), $shortrealtobits(4), $shortrealtobits(5), $shortrealtobits(1), $shortrealtobits(2), $shortrealtobits(1), $shortrealtobits(8), $shortrealtobits(2), $shortrealtobits(9), $shortrealtobits(3), $shortrealtobits(9), $shortrealtobits(3), $shortrealtobits(1), $shortrealtobits(3), $shortrealtobits(3), $shortrealtobits(7), $shortrealtobits(6), $shortrealtobits(2), $shortrealtobits(7), $shortrealtobits(2), $shortrealtobits(8), $shortrealtobits(10), $shortrealtobits(2), $shortrealtobits(2), $shortrealtobits(10), $shortrealtobits(10), $shortrealtobits(9), $shortrealtobits(9), $shortrealtobits(4), $shortrealtobits(3), $shortrealtobits(2), $shortrealtobits(9), $shortrealtobits(5), $shortrealtobits(4), $shortrealtobits(9), $shortrealtobits(2), $shortrealtobits(1), $shortrealtobits(6), $shortrealtobits(5), $shortrealtobits(4), $shortrealtobits(10), $shortrealtobits(6), $shortrealtobits(3), $shortrealtobits(6), $shortrealtobits(9), $shortrealtobits(9), $shortrealtobits(4), $shortrealtobits(7), $shortrealtobits(5), $shortrealtobits(2), $shortrealtobits(2), $shortrealtobits(7), $shortrealtobits(6), $shortrealtobits(3), $shortrealtobits(9), $shortrealtobits(9), $shortrealtobits(7), $shortrealtobits(2), $shortrealtobits(9), $shortrealtobits(1), $shortrealtobits(10), $shortrealtobits(7), $shortrealtobits(10), $shortrealtobits(1), $shortrealtobits(3), $shortrealtobits(9), $shortrealtobits(4), $shortrealtobits(4), $shortrealtobits(4), $shortrealtobits(6), $shortrealtobits(7), $shortrealtobits(5), $shortrealtobits(5), $shortrealtobits(6), $shortrealtobits(3), $shortrealtobits(5), $shortrealtobits(4), $shortrealtobits(8), $shortrealtobits(8), $shortrealtobits(5), $shortrealtobits(3), $shortrealtobits(10), $shortrealtobits(6), $shortrealtobits(6), $shortrealtobits(8), $shortrealtobits(3), $shortrealtobits(8), $shortrealtobits(9), $shortrealtobits(7), $shortrealtobits(9), $shortrealtobits(4), $shortrealtobits(8), $shortrealtobits(2), $shortrealtobits(9), $shortrealtobits(2), $shortrealtobits(5), $shortrealtobits(9), $shortrealtobits(4), $shortrealtobits(8), $shortrealtobits(6), $shortrealtobits(8), $shortrealtobits(1), $shortrealtobits(6), $shortrealtobits(10), $shortrealtobits(5), $shortrealtobits(5), $shortrealtobits(4), $shortrealtobits(1), $shortrealtobits(8), $shortrealtobits(9), $shortrealtobits(10), $shortrealtobits(5), $shortrealtobits(10), $shortrealtobits(7), $shortrealtobits(9), $shortrealtobits(5), $shortrealtobits(8), $shortrealtobits(2), $shortrealtobits(3), $shortrealtobits(9), $shortrealtobits(4), $shortrealtobits(1), $shortrealtobits(3), $shortrealtobits(5), $shortrealtobits(9), $shortrealtobits(8), $shortrealtobits(4), $shortrealtobits(9), $shortrealtobits(1), $shortrealtobits(1), $shortrealtobits(10), $shortrealtobits(7), $shortrealtobits(9), $shortrealtobits(9), $shortrealtobits(9), $shortrealtobits(1), $shortrealtobits(8), $shortrealtobits(5)};

  always_ff @(posedge clock) begin
    if (read) readdata <= {mem[address+7], mem[address+6], mem[address+5], mem[address+4],
                       mem[address+3], mem[address+2], mem[address+1], mem[address]};
    else readdata <= 'b0;
  end

endmodule: fakemem_readA


module fakemem_readB
  (input logic read, clock, 
   input logic [`ADDR_WIDTH-1:0] address,
   output logic [`BANDWIDTH-1:0][`DATA_WIDTH-1:0] readdata);

  logic [511:0][31:0] mem;

  assign mem[383:0] = {$shortrealtobits(2), $shortrealtobits(4), $shortrealtobits(6), $shortrealtobits(2), $shortrealtobits(5), $shortrealtobits(5), $shortrealtobits(8), $shortrealtobits(7), $shortrealtobits(8), $shortrealtobits(5), $shortrealtobits(6), $shortrealtobits(6), $shortrealtobits(6), $shortrealtobits(1), $shortrealtobits(7), $shortrealtobits(6), $shortrealtobits(2), $shortrealtobits(9), $shortrealtobits(5), $shortrealtobits(7), $shortrealtobits(9), $shortrealtobits(7), $shortrealtobits(7), $shortrealtobits(10), $shortrealtobits(5), $shortrealtobits(10), $shortrealtobits(3), $shortrealtobits(9), $shortrealtobits(10), $shortrealtobits(4), $shortrealtobits(3), $shortrealtobits(4), $shortrealtobits(7), $shortrealtobits(5), $shortrealtobits(4), $shortrealtobits(10), $shortrealtobits(5), $shortrealtobits(8), $shortrealtobits(5), $shortrealtobits(10), $shortrealtobits(4), $shortrealtobits(8), $shortrealtobits(9), $shortrealtobits(8), $shortrealtobits(2), $shortrealtobits(1), $shortrealtobits(6), $shortrealtobits(3), $shortrealtobits(5), $shortrealtobits(5), $shortrealtobits(8), $shortrealtobits(10), $shortrealtobits(2), $shortrealtobits(8), $shortrealtobits(2), $shortrealtobits(10), $shortrealtobits(6), $shortrealtobits(10), $shortrealtobits(7), $shortrealtobits(7), $shortrealtobits(1), $shortrealtobits(10), $shortrealtobits(7), $shortrealtobits(9), $shortrealtobits(3), $shortrealtobits(6), $shortrealtobits(2), $shortrealtobits(4), $shortrealtobits(9), $shortrealtobits(5), $shortrealtobits(4), $shortrealtobits(1), $shortrealtobits(9), $shortrealtobits(5), $shortrealtobits(6), $shortrealtobits(2), $shortrealtobits(10), $shortrealtobits(8), $shortrealtobits(7), $shortrealtobits(8), $shortrealtobits(4), $shortrealtobits(4), $shortrealtobits(7), $shortrealtobits(9), $shortrealtobits(4), $shortrealtobits(5), $shortrealtobits(9), $shortrealtobits(3), $shortrealtobits(8), $shortrealtobits(6), $shortrealtobits(2), $shortrealtobits(10), $shortrealtobits(2), $shortrealtobits(6), $shortrealtobits(2), $shortrealtobits(7), $shortrealtobits(7), $shortrealtobits(6), $shortrealtobits(7), $shortrealtobits(4), $shortrealtobits(2), $shortrealtobits(6), $shortrealtobits(10), $shortrealtobits(3), $shortrealtobits(8), $shortrealtobits(1), $shortrealtobits(3), $shortrealtobits(5), $shortrealtobits(6), $shortrealtobits(9), $shortrealtobits(9), $shortrealtobits(10), $shortrealtobits(6), $shortrealtobits(1), $shortrealtobits(6), $shortrealtobits(7), $shortrealtobits(5), $shortrealtobits(7), $shortrealtobits(10), $shortrealtobits(4), $shortrealtobits(8), $shortrealtobits(8), $shortrealtobits(8), $shortrealtobits(8), $shortrealtobits(4), $shortrealtobits(2), $shortrealtobits(8), $shortrealtobits(5), $shortrealtobits(6), $shortrealtobits(10), $shortrealtobits(1), $shortrealtobits(2), $shortrealtobits(2), $shortrealtobits(4), $shortrealtobits(5), $shortrealtobits(4), $shortrealtobits(5), $shortrealtobits(5), $shortrealtobits(4), $shortrealtobits(2), $shortrealtobits(7), $shortrealtobits(1), $shortrealtobits(3), $shortrealtobits(4), $shortrealtobits(3), $shortrealtobits(8), $shortrealtobits(8), $shortrealtobits(1), $shortrealtobits(5), $shortrealtobits(2), $shortrealtobits(1), $shortrealtobits(8), $shortrealtobits(5), $shortrealtobits(4), $shortrealtobits(4), $shortrealtobits(10), $shortrealtobits(1), $shortrealtobits(6), $shortrealtobits(7), $shortrealtobits(1), $shortrealtobits(8), $shortrealtobits(7), $shortrealtobits(2), $shortrealtobits(3), $shortrealtobits(3), $shortrealtobits(4), $shortrealtobits(6), $shortrealtobits(10), $shortrealtobits(5), $shortrealtobits(8), $shortrealtobits(6), $shortrealtobits(5), $shortrealtobits(10), $shortrealtobits(6), $shortrealtobits(6), $shortrealtobits(3), $shortrealtobits(8), $shortrealtobits(5), $shortrealtobits(1), $shortrealtobits(6), $shortrealtobits(9), $shortrealtobits(2), $shortrealtobits(1), $shortrealtobits(3), $shortrealtobits(4), $shortrealtobits(3), $shortrealtobits(7), $shortrealtobits(3), $shortrealtobits(7), $shortrealtobits(1), $shortrealtobits(10), $shortrealtobits(3), $shortrealtobits(9), $shortrealtobits(6), $shortrealtobits(8), $shortrealtobits(9), $shortrealtobits(10), $shortrealtobits(7), $shortrealtobits(7), $shortrealtobits(7), $shortrealtobits(9), $shortrealtobits(10), $shortrealtobits(4), $shortrealtobits(10), $shortrealtobits(8), $shortrealtobits(5), $shortrealtobits(10), $shortrealtobits(5), $shortrealtobits(1), $shortrealtobits(4), $shortrealtobits(3), $shortrealtobits(3), $shortrealtobits(2), $shortrealtobits(2), $shortrealtobits(10), $shortrealtobits(8), $shortrealtobits(7), $shortrealtobits(8), $shortrealtobits(6), $shortrealtobits(6), $shortrealtobits(5), $shortrealtobits(9), $shortrealtobits(3), $shortrealtobits(3), $shortrealtobits(8), $shortrealtobits(9), $shortrealtobits(6), $shortrealtobits(7), $shortrealtobits(8), $shortrealtobits(4), $shortrealtobits(5), $shortrealtobits(1), $shortrealtobits(7), $shortrealtobits(7), $shortrealtobits(8), $shortrealtobits(9), $shortrealtobits(3), $shortrealtobits(5), $shortrealtobits(6), $shortrealtobits(7), $shortrealtobits(6), $shortrealtobits(7), $shortrealtobits(9), $shortrealtobits(6), $shortrealtobits(1), $shortrealtobits(8), $shortrealtobits(2), $shortrealtobits(5), $shortrealtobits(7), $shortrealtobits(8), $shortrealtobits(9), $shortrealtobits(10), $shortrealtobits(4), $shortrealtobits(9), $shortrealtobits(1), $shortrealtobits(4), $shortrealtobits(7), $shortrealtobits(8), $shortrealtobits(3), $shortrealtobits(3), $shortrealtobits(2), $shortrealtobits(9), $shortrealtobits(6), $shortrealtobits(5), $shortrealtobits(8), $shortrealtobits(3), $shortrealtobits(4), $shortrealtobits(6), $shortrealtobits(7), $shortrealtobits(6), $shortrealtobits(10), $shortrealtobits(7), $shortrealtobits(7), $shortrealtobits(10), $shortrealtobits(1), $shortrealtobits(9), $shortrealtobits(10), $shortrealtobits(5), $shortrealtobits(7), $shortrealtobits(4), $shortrealtobits(1), $shortrealtobits(1), $shortrealtobits(5), $shortrealtobits(7), $shortrealtobits(7), $shortrealtobits(8), $shortrealtobits(4), $shortrealtobits(8), $shortrealtobits(4), $shortrealtobits(3), $shortrealtobits(10), $shortrealtobits(4), $shortrealtobits(8), $shortrealtobits(9), $shortrealtobits(9), $shortrealtobits(4), $shortrealtobits(4), $shortrealtobits(8), $shortrealtobits(4), $shortrealtobits(7), $shortrealtobits(8), $shortrealtobits(10), $shortrealtobits(9), $shortrealtobits(6), $shortrealtobits(4), $shortrealtobits(8), $shortrealtobits(1), $shortrealtobits(4), $shortrealtobits(1), $shortrealtobits(2), $shortrealtobits(5), $shortrealtobits(8), $shortrealtobits(9), $shortrealtobits(1), $shortrealtobits(3), $shortrealtobits(5), $shortrealtobits(9), $shortrealtobits(9), $shortrealtobits(9), $shortrealtobits(10), $shortrealtobits(2), $shortrealtobits(4), $shortrealtobits(3), $shortrealtobits(8), $shortrealtobits(7), $shortrealtobits(9), $shortrealtobits(1), $shortrealtobits(4), $shortrealtobits(6), $shortrealtobits(1), $shortrealtobits(4), $shortrealtobits(9), $shortrealtobits(6), $shortrealtobits(7), $shortrealtobits(1), $shortrealtobits(7), $shortrealtobits(6), $shortrealtobits(6), $shortrealtobits(10), $shortrealtobits(5), $shortrealtobits(2), $shortrealtobits(5), $shortrealtobits(8), $shortrealtobits(9), $shortrealtobits(8), $shortrealtobits(1), $shortrealtobits(7), $shortrealtobits(10), $shortrealtobits(10), $shortrealtobits(10), $shortrealtobits(8), $shortrealtobits(1), $shortrealtobits(6), $shortrealtobits(2), $shortrealtobits(10), $shortrealtobits(4), $shortrealtobits(4), $shortrealtobits(3), $shortrealtobits(3), $shortrealtobits(8), $shortrealtobits(4), $shortrealtobits(3), $shortrealtobits(3), $shortrealtobits(8), $shortrealtobits(7), $shortrealtobits(1), $shortrealtobits(5), $shortrealtobits(4), $shortrealtobits(1), $shortrealtobits(10), $shortrealtobits(7), $shortrealtobits(4), $shortrealtobits(9), $shortrealtobits(3), $shortrealtobits(1), $shortrealtobits(7), $shortrealtobits(2), $shortrealtobits(9), $shortrealtobits(1), $shortrealtobits(4), $shortrealtobits(8), $shortrealtobits(2), $shortrealtobits(9), $shortrealtobits(7)};

  always_ff @(posedge clock) begin
    if (read) readdata <= {mem[address+7], mem[address+6], mem[address+5], mem[address+4],
                       mem[address+3], mem[address+2], mem[address+1], mem[address]};
    else readdata <= 'b0;
  end

endmodule: fakemem_readB


module fakemem_write
  (input logic write, clock, 
   input logic [`ADDR_WIDTH-1:0] address,
   input logic [`BANDWIDTH-1:0][`DATA_WIDTH-1:0] writedata);

  logic [511:0][31:0] mem;

  always_ff @(posedge clock) begin
    if (write) {mem[address+7], mem[address+6], mem[address+5], mem[address+4],
                mem[address+3], mem[address+2], mem[address+1], mem[address]} <= writedata;
  end

endmodule: fakemem_write


module fakemem
  (input logic read, write, clock, 
   input logic [`ADDR_WIDTH-1:0] address,
   input logic [`DATA_WIDTH*`BANDWIDTH-1:0] writedata,
   output logic [`DATA_WIDTH*`BANDWIDTH-1:0] readdata);

  logic [63:0][255:0] mem;

  always_comb begin
    mem[0] = {MAT_SCAL_MUL, 14'd128, 7'd8, 7'd16};
    mem[1] = $shortrealtobits(3);
  end

  always_ff @(posedge clock) begin
    if (read) readdata <= mem[address];
    // else if (write) mem[address] <= writedata;
    else readdata <= 'b0;
  end

endmodule: fakemem