`define SIZE_MAX 128

`define OP_ADDR 0
`define SCALAR_ADDR 1
`define DATAA_ADDR 10
`define DATAB_ADDR 30
`define RES_ADDR 50

`define ADDR_WIDTH 14
`define DATA_WIDTH 32
`define OP_WIDTH 4
`define DIM_WIDTH 7

`define BANDWIDTH 4

`define SINGLE_ACCESS 8

`define CYCLE_WIDTH 4
`define CYCLE_MUL 5
`define CYCLE_DIV 5
`define CYCLE_ADD 7
`define CYCLE_INV 5
`define CYCLE_MAT_MUL 5

`timescale 1 ps / 1 ps